module decoder5to32(input [4:0] offset, output reg [31:0] outputReg);
	always @(offset)
	begin
		case(offset)
			5'd0  : outputReg = 32'b00000000000000000000000000000001;
			5'd1  : outputReg = 32'b00000000000000000000000000000010;
			5'd2  : outputReg = 32'b00000000000000000000000000000100;
			5'd3  : outputReg = 32'b00000000000000000000000000001000;
			5'd4  : outputReg = 32'b00000000000000000000000000010000;
			5'd5  : outputReg = 32'b00000000000000000000000000100000;
			5'd6  : outputReg = 32'b00000000000000000000000001000000;
			5'd7  : outputReg = 32'b00000000000000000000000010000000;
			5'd8  : outputReg = 32'b00000000000000000000000100000000;
			5'd9  : outputReg = 32'b00000000000000000000001000000000;
			5'd10 : outputReg = 32'b00000000000000000000010000000000;
			5'd11 : outputReg = 32'b00000000000000000000100000000000;
			5'd12 : outputReg = 32'b00000000000000000001000000000000;
			5'd13 : outputReg = 32'b00000000000000000010000000000000;
			5'd14 : outputReg = 32'b00000000000000000100000000000000;
			5'd15 : outputReg = 32'b00000000000000001000000000000000;
			5'd16 : outputReg = 32'b00000000000000010000000000000000;
			5'd17 : outputReg = 32'b00000000000000100000000000000000;
			5'd18 : outputReg = 32'b00000000000001000000000000000000;
			5'd19 : outputReg = 32'b00000000000010000000000000000000;
			5'd20 : outputReg = 32'b00000000000100000000000000000000;
			5'd21 : outputReg = 32'b00000000001000000000000000000000;
			5'd22 : outputReg = 32'b00000000010000000000000000000000;
			5'd23 : outputReg = 32'b00000000100000000000000000000000;
			5'd24 : outputReg = 32'b00000001000000000000000000000000;
			5'd25 : outputReg = 32'b00000010000000000000000000000000;
			5'd26 : outputReg = 32'b00000100000000000000000000000000;
			5'd27 : outputReg = 32'b00001000000000000000000000000000;
			5'd28 : outputReg = 32'b00010000000000000000000000000000;
			5'd29 : outputReg = 32'b00100000000000000000000000000000;
			5'd30 : outputReg = 32'b01000000000000000000000000000000;
			5'd31 : outputReg = 32'b10000000000000000000000000000000;
		endcase
	end
endmodule