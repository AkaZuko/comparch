module register32bit_normal(input clk, input reset, input regWrite, input decOut1b, input [31:0] writeData, output  [31:0] outR );
	D_ff_normal d0(clk, reset, regWrite, decOut1b, writeData[0], outR[0]);
	D_ff_normal d1(clk, reset, regWrite, decOut1b, writeData[1], outR[1]);
	D_ff_normal d2(clk, reset, regWrite, decOut1b, writeData[2], outR[2]);
	D_ff_normal d3(clk, reset, regWrite, decOut1b, writeData[3], outR[3]);
	D_ff_normal d4(clk, reset, regWrite, decOut1b, writeData[4], outR[4]);
	D_ff_normal d5(clk, reset, regWrite, decOut1b, writeData[5], outR[5]);
	D_ff_normal d6(clk, reset, regWrite, decOut1b, writeData[6], outR[6]);
	D_ff_normal d7(clk, reset, regWrite, decOut1b, writeData[7], outR[7]);
	D_ff_normal d8(clk, reset, regWrite, decOut1b, writeData[8], outR[8]);
	D_ff_normal d9(clk, reset, regWrite, decOut1b, writeData[9], outR[9]);
	D_ff_normal d10(clk, reset, regWrite, decOut1b, writeData[10], outR[10]);
	D_ff_normal d11(clk, reset, regWrite, decOut1b, writeData[11], outR[11]);
	D_ff_normal d12(clk, reset, regWrite, decOut1b, writeData[12], outR[12]);
	D_ff_normal d13(clk, reset, regWrite, decOut1b, writeData[13], outR[13]);
	D_ff_normal d14(clk, reset, regWrite, decOut1b, writeData[14], outR[14]);
	D_ff_normal d15(clk, reset, regWrite, decOut1b, writeData[15], outR[15]);

	D_ff_normal d16(clk, reset, regWrite, decOut1b, writeData[16], outR[16]);
	D_ff_normal d17(clk, reset, regWrite, decOut1b, writeData[17], outR[17]);
	D_ff_normal d18(clk, reset, regWrite, decOut1b, writeData[18], outR[18]);
	D_ff_normal d19(clk, reset, regWrite, decOut1b, writeData[19], outR[19]);
	D_ff_normal d20(clk, reset, regWrite, decOut1b, writeData[20], outR[20]);
	D_ff_normal d21(clk, reset, regWrite, decOut1b, writeData[21], outR[21]);
	D_ff_normal d22(clk, reset, regWrite, decOut1b, writeData[22], outR[22]);
	D_ff_normal d23(clk, reset, regWrite, decOut1b, writeData[23], outR[23]);
	D_ff_normal d24(clk, reset, regWrite, decOut1b, writeData[24], outR[24]);
	D_ff_normal d25(clk, reset, regWrite, decOut1b, writeData[25], outR[25]);
	D_ff_normal d26(clk, reset, regWrite, decOut1b, writeData[26], outR[26]);
	D_ff_normal d27(clk, reset, regWrite, decOut1b, writeData[27], outR[27]);
	D_ff_normal d28(clk, reset, regWrite, decOut1b, writeData[28], outR[28]);
	D_ff_normal d29(clk, reset, regWrite, decOut1b, writeData[29], outR[29]);
	D_ff_normal d30(clk, reset, regWrite, decOut1b, writeData[30], outR[30]);
	D_ff_normal d31(clk, reset, regWrite, decOut1b, writeData[31], outR[31]);
endmodule