module IFID(input clk, input reset, input IFwrite, input IFflush,)